--blank 
